
----------------------------------------------------------------
-- Instruction Memory
----------------------------------------------------------------
constant INSTR_MEM : MEM_128x32 := (		x"E59F11F8", 
											x"E59F21F8", 
											x"E59F3200", 
											x"E5924000", 
											x"E5814000", 
											x"E2533001", 
											x"1AFFFFFD", 
											x"E3530000", 
											x"0AFFFFF8", 
											x"EAFFFFFE", 
											others => x"00000000");

----------------------------------------------------------------
-- Data (Constant) Memory
----------------------------------------------------------------
constant DATA_CONST_MEM : MEM_128x32 := (	x"00000C00", 
											x"00000C04", 
											x"00000C08", 
											x"00000C0C", 
											x"00000004", 
											x"00000800", 
											x"ABCD1234", 
											x"6C6C6548", 
											x"6F57206F", 
											x"21646C72", 
											x"00212121", 
											others => x"00000000");

